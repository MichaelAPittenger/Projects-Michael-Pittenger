LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Problem_4_48 IS
	PORT(	X1, X2, X3, X4	: IN	STD_LOGIC;
			f					: OUT	STD_LOGIC);
END Problem_4_48;

ARCHITECTURE Structure OF Problem_4_48 IS

BEGIN

	f <= (NOT X1 AND NOT X2 AND NOT X4) OR 
		  (NOT X1 AND NOT X3) OR 
		  (NOT X1 AND X2 AND X4) OR 
		  (NOT X2 AND NOT X3) OR 
		  (X1 AND X3 AND X4) OR 
		  (X1 AND X2 AND NOT X4);

END Structure;