LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Project1 IS
	PORT(	SW			: IN  STD_LOGIC_VECTOR(9 DOWNTO 0);
			KEY		: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
			LEDR		: OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
			CLOCK_50	: IN STD_LOGIC;
			HEX0		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX1		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX2		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX3		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX4		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX5		: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END Project1;

ARCHITECTURE Structure OF Project1 IS

	--Components
	COMPONENT adder4
		PORT (	Cin    : IN    STD_LOGIC;
					X, Y   : IN    STD_LOGIC_VECTOR(3 DOWNTO 0);
					S      : OUT   STD_LOGIC_VECTOR(3 DOWNTO 0);
					Cout   : OUT   STD_LOGIC);
	END COMPONENT;
	
	COMPONENT MUX_12TO4 
		PORT(	S		: IN	STD_LOGIC_VECTOR(1 DOWNTO 0);
				A, B, C	: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
				Y			: OUT	STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT MUX_8TO4 IS
		PORT(	S		: IN	STD_LOGIC;
				A, B	: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
				Y		: OUT	STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT BCD IS
		PORT(	I				: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
				Out1, Out0	: OUT	STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT sevenSeg IS
		PORT(	d0		: IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
				HEX	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0));
	END COMPONENT;
	
	--Signals
	SIGNAL A, B, nB, C, ZERO, MUX3TO1, MUX2TO1, SUM, AXORB	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL Cin, Cout, C3, C2, C1, S1, S0				:	STD_LOGIC;
	SIGNAL D5, D4, D3, D2, D1, D0							:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	
BEGIN

	--DFF INPUT
	PROCESS(CLOCK_50)
	BEGIN
		IF CLOCK_50'EVENT AND CLOCK_50 ='1' THEN
			A <= SW(7 DOWNTO 4);
			B <= SW(3 DOWNTO 0);
			S1 <= SW(9);
			S0 <= SW(8);	
			Cin <= NOT KEY(0);
		END IF;
	END PROCESS;
	
	--DFF OUTPUT
	PROCESS(CLOCK_50)
	BEGIN
		IF CLOCK_50'EVENT AND CLOCK_50 ='0' THEN
			C <= MUX2TO1;
		END IF;
	END PROCESS;

	--OTHER SIGNALS
	nB <= NOT B;
	ZERO <= "0000";
	
	C3 <= NOT S1 OR NOT S0;
	C2 <= NOT S1 AND NOT S0;
	C1 <= S1 AND NOT S0;

	--MUX TEST
	LEDR(9 DOWNTO 4) <= "000000";
	
	--12TO4 MUX - 2 SEL BITS
	MICHAEL0	: MUX_12TO4 PORT MAP ((C2 & C1), B, nB, ZERO, MUX3TO1);
	
	--4-BIT ADDER
	MICHAEL1	: adder4 PORT MAP(Cin, A, MUX3TO1, SUM, Cout);
	
	--XOR
	AXORB <= A XOR B;
	
	--8TO4 MUX - 1 SEL BIT
	MICHAEL2	: MUX_8TO4 PORT MAP (C3, SUM, AXORB, MUX2TO1);
	
	--LED OUTPUT
	LEDR(3 DOWNTO 0) <= C;
	

	--SEVEN SEGMENT DISPLAY
	MICHAEL3	: BCD PORT MAP (A, D5, D4);
	MICHAEL4	: BCD PORT MAP (B, D3, D2);
	MICHAEL5	: BCD PORT MAP (C, D1, D0);
	
	MICHAEL6		: sevenSeg PORT MAP (D5, HEX5);
	MICHAEL7		: sevenSeg PORT MAP (D4, HEX4);
	MICHAEL8		: sevenSeg PORT MAP (D3, HEX3);
	MICHAEL9		: sevenSeg PORT MAP (D2, HEX2);
	MICHAEL10	: sevenSeg PORT MAP (D1, HEX1);
	MICHAEL11	: sevenSeg PORT MAP (D0, HEX0);
	

END Structure;