LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PROBLEM_7_10 IS
	PORT(	CLK	: IN	STD_LOGIC;
			CLR	: IN	STD_LOGIC;
			T		: IN	STD_LOGIC;
			Q		: OUT	STD_LOGIC;
			nQ		: OUT	STD_LOGIC);
END PROBLEM_7_10;

ARCHITECTURE BEHAVIORAL OF PROBLEM_7_10 IS

		SIGNAL Q_INT : STD_LOGIC := '0';

BEGIN

	PROCESS(CLK, CLR)
	BEGIN
		IF CLR = '1' THEN
			Q_INT <= '0';
		ELSIF CLK'EVENT AND CLK = '1' THEN
			IF T = '1' THEN
				Q_INT <= NOT Q_INT;
			END IF;
		END IF;
	END PROCESS;
	
	Q <= Q_INT;

END BEHAVIORAL;