LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Problem_4_49 IS
	PORT(	X1, X2, X3, X4	: IN	STD_LOGIC;
			f					: OUT	STD_LOGIC);
END Problem_4_49;

ARCHITECTURE Structure OF Problem_4_49 IS

BEGIN

	f <= (NOT X1 AND NOT X3) OR 
		  (X1 AND X2 AND X3) OR 
		  (NOT X1 AND X2 AND X4);

END Structure;