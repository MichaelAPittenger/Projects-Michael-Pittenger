--Michael Pittenger
--EE 421/621

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY VHDLHW IS
    PORT(	SW		: IN  STD_LOGIC_VECTOR(7 DOWNTO 0);
				LEDR	: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
				HEX0	: OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
				HEX1	: OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END VHDLHW;

ARCHITECTURE LogicFunc OF VHDLHW IS

	--Components
	COMPONENT adder4
		PORT (	Cin    : IN    STD_LOGIC;
					X, Y   : IN    STD_LOGIC_VECTOR(3 DOWNTO 0);
					S      : OUT   STD_LOGIC_VECTOR(3 DOWNTO 0);
					Cout   : OUT   STD_LOGIC);
	END COMPONENT;
	
	COMPONENT sevenSeg
		PORT(	d0		: IN 	STD_LOGIC_VECTOR(3 DOWNTO 0);
				HEX	: OUT	STD_LOGIC_VECTOR(6 DOWNTO 0));	
	END COMPONENT;
	
	COMPONENT BCD
		PORT(	I				: IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
				Out1, Out0	: OUT	STD_LOGIC_VECTOR(3 DOWNTO 0));
	END COMPONENT;

	--Signals
	SIGNAL Cin 	: STD_LOGIC := '0';
	SIGNAL Cout	: STD_LOGIC;
	SIGNAL S		: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL d0 	: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL d1 	: STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN

	--4-bit Adder
	michael: adder4 PORT MAP (Cin, SW(7 DOWNTO 4), SW(3 DOWNTO 0), S(3 DOWNTO 0), Cout);

	--Binary Coded Decimal
	michael0: BCD PORT MAP (S(3 DOWNTO 0), d1(3 DOWNTO 0), d0(3 DOWNTO 0));
	
	--Seven Segment Display[
	michael1: sevenSeg PORT MAP (d0(3 DOWNTO 0), HEX0(6 DOWNTO 0));
	michael2: sevenSeg PORT MAP (d1(3 DOWNTO 0), HEX1(6 DOWNTO 0));

END LogicFunc;
