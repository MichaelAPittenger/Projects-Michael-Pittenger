LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY Problem_4_46 IS
	PORT(	X1, X2, X3, X4, X5, X6, X7	: IN	STD_LOGIC;
			f									: OUT	STD_LOGIC);
END Problem_4_46;

ARCHITECTURE Structure OF Problem_4_46 IS

	SIGNAL W1, W23, W123, W5, W6, W7, W56, W456, W4567, W1234567	: STD_LOGIC;

BEGIN

	W1			<= NOT (X1 AND X1);
	W23		<= NOT (X2 AND X3);
	W123		<= NOT (W1 AND W23);
	
	W5			<= NOT (X5 AND X5);
	W6			<= NOT (X6 AND X6);
	W56		<= NOT (W5 AND W6);
	W456		<= NOT (X4 AND W56);
	
	W7			<= NOT (X7 AND X7);
	W4567		<= NOT (W456 AND W7);
	W1234567	<= NOT (W123 AND W4567);
	
	f			<= NOT (W1234567 AND W1234567);

END Structure;