LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY PROBLEM_7_23 IS
	PORT(	clk		: IN	STD_LOGIC;
			reset		: IN	STD_LOGIC;
			Q			: OUT	STD_LOGIC_VECTOR(3 DOWNTO 0));
END PROBLEM_7_23;

ARCHITECTURE BEHAVIORAL OF PROBLEM_7_23 IS

	SIGNAL count : STD_LOGIC_VECTOR(3 DOWNTO 0) := '0000';

BEGIN

	PROCESS (clk)
	BEGIN
		IF RISING_EDGE(clk) THEN
			IF reset = '1' THEN
				count <= '0000';
			ELSIF count <= '1011' THEN
				count <= '0000';
			ELSE
				count <= count + 1;
		END IF;
	END PROCESS;
	
	Q <= count;

END BEHAVIORAL;
